.subckt ORG_CAVLC_COMPLEX4_06W GND cl3#A cl1#B VCC cl0#Y cl2#B cl2#Y cl2#A cl3#C cl3#B cl1#Y cl1#A
Mcl0#0 cl0#a_9_54# cl1#Y VCC VCC PMOS_VTL W=0.6u L=0.05u
+ ad=0p pd=0u as=0p ps=0u 
Mcl0#1 cl0#Y cl2#Y cl0#a_9_54# VCC PMOS_VTL W=0.6u L=0.05u
+ ad=0p pd=0u as=0p ps=0u 
Mcl0#2 VCC cl3#Y cl0#Y VCC PMOS_VTL W=0.3u L=0.05u
+ ad=0p pd=0u as=0p ps=0u 
Mcl0#3 GND cl1#Y cl0#a_2_6# GND NMOS_VTL W=0.3u L=0.05u
+ ad=0p pd=0u as=0p ps=0u 
Mcl0#4 cl0#a_2_6# cl2#Y GND GND NMOS_VTL W=0.3u L=0.05u
+ ad=0p pd=0u as=0p ps=0u 
Mcl0#5 cl0#Y cl3#Y cl0#a_2_6# GND NMOS_VTL W=0.3u L=0.05u
+ ad=0p pd=0u as=0p ps=0u 
Mcl1#0 cl1#Y cl1#A VCC VCC PMOS_VTL W=0.3u L=0.05u
+ ad=0p pd=0u as=0p ps=0u 
Mcl1#1 VCC cl1#B cl1#Y VCC PMOS_VTL W=0.3u L=0.05u
+ ad=0p pd=0u as=0p ps=0u 
Mcl1#2 cl1#a_9_6# cl1#A GND GND NMOS_VTL W=0.3u L=0.05u
+ ad=0p pd=0u as=0p ps=0u 
Mcl1#3 cl1#Y cl1#B cl1#a_9_6# GND NMOS_VTL W=0.3u L=0.05u
+ ad=0p pd=0u as=0p ps=0u 
Mcl2#0 cl2#Y cl2#A VCC VCC PMOS_VTL W=0.3u L=0.05u
+ ad=0p pd=0u as=0p ps=0u 
Mcl2#1 VCC cl2#B cl2#Y VCC PMOS_VTL W=0.3u L=0.05u
+ ad=0p pd=0u as=0p ps=0u 
Mcl2#2 cl2#a_9_6# cl2#A GND GND NMOS_VTL W=0.3u L=0.05u
+ ad=0p pd=0u as=0p ps=0u 
Mcl2#3 cl2#Y cl2#B cl2#a_9_6# GND NMOS_VTL W=0.3u L=0.05u
+ ad=0p pd=0u as=0p ps=0u 
Mcl3#0 cl3#Y cl3#A VCC VCC PMOS_VTL W=0.3u L=0.05u
+ ad=0p pd=0u as=0p ps=0u 
Mcl3#1 VCC cl3#B cl3#Y VCC PMOS_VTL W=0.3u L=0.05u
+ ad=0p pd=0u as=0p ps=0u 
Mcl3#2 cl3#Y cl3#C VCC VCC PMOS_VTL W=0.3u L=0.05u
+ ad=0p pd=0u as=0p ps=0u 
Mcl3#3 cl3#a_9_6# cl3#A GND GND NMOS_VTL W=0.45u L=0.05u
+ ad=0p pd=0u as=0p ps=0u 
Mcl3#4 cl3#a_14_6# cl3#B cl3#a_9_6# GND NMOS_VTL W=0.45u L=0.05u
+ ad=0p pd=0u as=0p ps=0u 
Mcl3#5 cl3#Y cl3#C cl3#a_14_6# GND NMOS_VTL W=0.45u L=0.05u
+ ad=0p pd=0u as=0p ps=0u 
.ends ORG_CAVLC_COMPLEX4_06W
* pattern code: [OAI21X1,NAND2X1,NAND2X1,NAND3X1]
* 5 occurrences in design 
* each contains 4 cells
* Example occurence:
*   .subckt OAI21X1 A=$abc$3639$new_n126_ B=$abc$3639$new_n135_ C=$abc$3639$new_n141_ Y=$abc$3639$new_n142_
*   .subckt NAND2X1 A=ctable[0] B=$abc$3639$new_n30_ Y=$abc$3639$new_n126_
*   .subckt NAND2X1 A=trailingones[1] B=$abc$3639$new_n27_ Y=$abc$3639$new_n135_
*   .subckt NAND3X1 A=totalcoeffs[0] B=$abc$3639$new_n139_ C=$abc$3639$new_n140_ Y=$abc$3639$new_n141_

.subckt BAR_COMPLEX1_06W GND VCC Y a b c d e f g h i j k 
M0 Y i pN4 VCC PMOS_VTL W=0.6u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M1 pN2 b pN1 VCC PMOS_VTL W=1.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M2 pN2 a pN1 VCC PMOS_VTL W=1.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M3 Y c pN3 VCC PMOS_VTL W=1.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M4 pN1 e pN4 VCC PMOS_VTL W=1.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M5 pN1 f pN4 VCC PMOS_VTL W=1.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M6 pN3 g pN2 VCC PMOS_VTL W=1.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M7 pN3 h pN2 VCC PMOS_VTL W=1.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M8 Y d pN3 VCC PMOS_VTL W=1.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M9 pN4 j VCC VCC PMOS_VTL W=1.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M10 pN4 k VCC VCC PMOS_VTL W=1.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M11 nN1 k GND GND NMOS_VTL W=0.3u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M12 nN2 b nN3 GND NMOS_VTL W=0.45u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M13 Y a nN2 GND NMOS_VTL W=0.45u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M14 nN4 d nN3 GND NMOS_VTL W=0.45u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M15 nN5 e nN3 GND NMOS_VTL W=0.45u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M16 Y c nN4 GND NMOS_VTL W=0.45u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M17 Y f nN5 GND NMOS_VTL W=0.45u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M18 nN6 h nN3 GND NMOS_VTL W=0.45u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M19 nN3 i GND GND NMOS_VTL W=0.45u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M20 Y g nN6 GND NMOS_VTL W=0.45u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M21 Y j nN1 GND NMOS_VTL W=0.3u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
.ends BAR_COMPLEX1_06W

.subckt LOG2_COMPLEX6_06W GND VCC Y a b c d e f 
M0 Y INVY VCC VCC PMOS W=0.3u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M1 pN2 b pN1 VCC PMOS W=0.9u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M2 INVY c pN2 VCC PMOS W=0.9u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M3 INVY d pN2 VCC PMOS W=0.9u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M4 pN1 e VCC VCC PMOS W=0.9u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M5 pN1 f VCC VCC PMOS W=0.9u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M6 pN2 a pN1 VCC PMOS W=0.9u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M7 nN1 a GND GND NMOS W=0.3u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M8 INVY b nN1 GND NMOS W=0.3u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M9 nN3 c GND GND NMOS W=0.3u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M10 INVY d nN3 GND NMOS W=0.3u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M11 INVY e nN2 GND NMOS W=0.3u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M12 nN2 f GND GND NMOS W=0.3u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M13 Y INVY GND GND NMOS W=0.15u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
.ends LOG2_COMPLEX6_06W

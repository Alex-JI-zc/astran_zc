.subckt COMPLEX7 GND VCC Y a b c 
M0 Y b pN2 VCC PMOS_VTL W=1.2u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M1 pN1 a VCC VCC PMOS_VTL W=1.2u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M2 pN2 c pN1 VCC PMOS_VTL W=1.2u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M3 Y c GND GND NMOS_VTL W=0.2u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M4 Y a GND GND NMOS_VTL W=0.2u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M5 Y b GND GND NMOS_VTL W=0.2u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
.ends COMPLEX7

.subckt COMPLEX101 GND VCC Y a b c d 
M0 Y INVY VCC VCC PMOS_VTL W=0.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M1 pN2 b pN1 VCC PMOS_VTL W=1.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M2 pN1 c VCC VCC PMOS_VTL W=1.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M3 INVY d VCC VCC PMOS_VTL W=0.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M4 INVY a pN2 VCC PMOS_VTL W=1.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M5 INVY a nN1 GND NMOS_VTL W=0.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M6 INVY b nN1 GND NMOS_VTL W=0.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M7 INVY c nN1 GND NMOS_VTL W=0.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M8 nN1 d GND GND NMOS_VTL W=0.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M9 Y INVY GND GND NMOS_VTL W=0.25u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
.ends COMPLEX101

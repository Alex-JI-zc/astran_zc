.subckt COMPLEX106 GND VCC Y a b c d e f g 
M0 Y INVY VCC VCC PMOS_VTL W=0.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M1 INVY b pN2 VCC PMOS_VTL W=1.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M2 pN1 c VCC VCC PMOS_VTL W=1.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M3 INVY d pN4 VCC PMOS_VTL W=1.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M4 pN4 e pN3 VCC PMOS_VTL W=1.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M5 pN3 f VCC VCC PMOS_VTL W=1.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M6 pN4 g VCC VCC PMOS_VTL W=1u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M7 pN2 a pN1 VCC PMOS_VTL W=1.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M8 INVY a nN2 GND NMOS_VTL W=0.75u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M9 INVY b nN2 GND NMOS_VTL W=0.75u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M10 INVY c nN2 GND NMOS_VTL W=0.75u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M11 nN2 d GND GND NMOS_VTL W=0.5u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M12 nN1 e GND GND NMOS_VTL W=0.75u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M13 nN1 f GND GND NMOS_VTL W=0.75u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M14 nN2 g nN1 GND NMOS_VTL W=0.75u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
M15 Y INVY GND GND NMOS_VTL W=0.25u L=0.05u 
+ ad=0p pd=0u as=0p ps=0u
.ends COMPLEX106
